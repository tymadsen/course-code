library ieee;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;
entity mod_n_counter is
	generic(
		N: natural;
		WIDTH: natural
	);
	port(
		clk, reset: in std_logic;
		en: in std_logic;
		q: out std_logic_vector (WIDTH-1 downto 0);
		pulse : out std_logic
	);
end mod_n_counter ;

architecture mod_arch of mod_n_counter is
	signal r_reg : unsigned (WIDTH-1 downto 0);
	signal r_next: unsigned(WIDTH-1 downto 0);
begin
	-- register
	process (clk, reset)
	begin
		if (reset ='1') then
			r_reg <= (others=>'0');
		elsif (clk'event and clk='1') then
			r_reg <= r_next;
		end if ;
	end process;
	-- next-state logic
	process (en, r_reg)
	begin
		r_next <= r_reg;
		if (en='1') then
			if r_reg=(N-1) then
				r_next <= (others=>'0');
			else
				r_next <= r_reg + 1;
			end if ;
		end if ;
	end process;
	-- output logic
	q <= std_logic_vector(r_reg);
	pulse <= '1' when r_reg=(N-1) else
	'0';
end mod_arch;